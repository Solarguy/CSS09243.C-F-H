module rom(out, address);
	output reg [63:0] out;
	input [7:0] address;
	
	always @(address) begin
		case (address)
			8'h00: out = 64'b0;
			8'h01: out = 64'b1;
			8'h02: out = 64'b10;
			8'h03: out = 64'b11;
			8'h04: out = 64'b100;
			8'h05: out = 64'b101;
			8'h06: out = 64'b110;
			8'h07: out = 64'b111;
			8'h08: out = 64'b1000;
			8'h09: out = 64'b1001;
			8'h0A: out = 64'b1010;
			8'h0B: out = 64'b1011;
			8'h0C: out = 64'b1100;
			8'h0D: out = 64'b1101;
			8'h0E: out = 64'b1110;
			8'h0F: out = 64'b1111;
			8'h10: out = 64'b10000;
			8'h11: out = 64'b10001;
			8'h12: out = 64'b10010;
			8'h13: out = 64'b10011;
			8'h14: out = 64'b10100;
			8'h15: out = 64'b10101;
			8'h16: out = 64'b10110;
			8'h17: out = 64'b10111;
			8'h18: out = 64'b11000;
			8'h19: out = 64'b11001;
			8'h1A: out = 64'b11010;
			8'h1B: out = 64'b11011;
			8'h1C: out = 64'b11100;
			8'h1D: out = 64'b11101;
			8'h1E: out = 64'b11110;
			8'h1F: out = 64'b11111;
			8'h20: out = 64'b100000;
			8'h21: out = 64'b100001;
			8'h22: out = 64'b100010;
			8'h23: out = 64'b100011;
			8'h24: out = 64'b100100;
			8'h25: out = 64'b100101;
			8'h26: out = 64'b100110;
			8'h27: out = 64'b100111;
			8'h28: out = 64'b101000;
			8'h29: out = 64'b101001;
			8'h2A: out = 64'b101010;
			8'h2B: out = 64'b101011;
			8'h2C: out = 64'b101100;
			8'h2D: out = 64'b101101;
			8'h2E: out = 64'b101110;
			8'h2F: out = 64'b101111;
			8'h30: out = 64'b110000;
			8'h31: out = 64'b110001;
			8'h32: out = 64'b110010;
			8'h33: out = 64'b110011;
			8'h34: out = 64'b110100;
			8'h35: out = 64'b110101;
			8'h36: out = 64'b110110;
			8'h37: out = 64'b110111;
			8'h38: out = 64'b111000;
			8'h39: out = 64'b111001;
			8'h3A: out = 64'b111010;
			8'h3B: out = 64'b111011;
			8'h3C: out = 64'b111100;
			8'h3D: out = 64'b111101;
			8'h3E: out = 64'b111110;
			8'h3F: out = 64'b111111;
			8'h40: out = 64'b0;
			8'h41: out = 64'b0;
			8'h42: out = 64'b0;
			8'h43: out = 64'b0;
			8'h44: out = 64'b0;
			8'h45: out = 64'b0;
			8'h46: out = 64'b0;
			8'h47: out = 64'b0;
			8'h48: out = 64'b0;
			8'h49: out = 64'b0;
			8'h4A: out = 64'b0;
			8'h4B: out = 64'b0;
			8'h4C: out = 64'b0;
			8'h4D: out = 64'b0;
			8'h4E: out = 64'b0;
			8'h4F: out = 64'b0;
			8'h50: out = 64'b0;
			8'h51: out = 64'b0;
			8'h52: out = 64'b0;
			8'h53: out = 64'b0;
			8'h54: out = 64'b0;
			8'h55: out = 64'b0;
			8'h56: out = 64'b0;
			8'h57: out = 64'b0;
			8'h58: out = 64'b0;
			8'h59: out = 64'b0;
			8'h5A: out = 64'b0;
			8'h5B: out = 64'b0;
			8'h5C: out = 64'b0;
			8'h5D: out = 64'b0;
			8'h5E: out = 64'b0;
			8'h5F: out = 64'b0;
			8'h60: out = 64'b0;
			8'h61: out = 64'b0;
			8'h62: out = 64'b0;
			8'h63: out = 64'b0;
			8'h64: out = 64'b0;
			8'h65: out = 64'b0;
			8'h66: out = 64'b0;
			8'h67: out = 64'b0;
			8'h68: out = 64'b0;
			8'h69: out = 64'b0;
			8'h6A: out = 64'b0;
			8'h6B: out = 64'b0;
			8'h6C: out = 64'b0;
			8'h6D: out = 64'b0;
			8'h6E: out = 64'b0;
			8'h6F: out = 64'b0;
			8'h70: out = 64'b0;
			8'h71: out = 64'b0;
			8'h72: out = 64'b0;
			8'h73: out = 64'b0;
			8'h74: out = 64'b0;
			8'h75: out = 64'b0;
			8'h76: out = 64'b0;
			8'h77: out = 64'b0;
			8'h78: out = 64'b0;
			8'h79: out = 64'b0;
			8'h7A: out = 64'b0;
			8'h7B: out = 64'b0;
			8'h7C: out = 64'b0;
			8'h7D: out = 64'b0;
			8'h7E: out = 64'b0;
			8'h7F: out = 64'b0;
			8'h80: out = 64'b0;
			8'h81: out = 64'b0;
			8'h82: out = 64'b0;
			8'h83: out = 64'b0;
			8'h84: out = 64'b0;
			8'h85: out = 64'b0;
			8'h86: out = 64'b0;
			8'h87: out = 64'b0;
			8'h88: out = 64'b0;
			8'h89: out = 64'b0;
			8'h8A: out = 64'b0;
			8'h8B: out = 64'b0;
			8'h8C: out = 64'b0;
			8'h8D: out = 64'b0;
			8'h8E: out = 64'b0;
			8'h8F: out = 64'b0;
			8'h90: out = 64'b0;
			8'h91: out = 64'b0;
			8'h92: out = 64'b0;
			8'h93: out = 64'b0;
			8'h94: out = 64'b0;
			8'h95: out = 64'b0;
			8'h96: out = 64'b0;
			8'h97: out = 64'b0;
			8'h98: out = 64'b0;
			8'h99: out = 64'b0;
			8'h9A: out = 64'b0;
			8'h9B: out = 64'b0;
			8'h9C: out = 64'b0;
			8'h9D: out = 64'b0;
			8'h9E: out = 64'b0;
			8'h9F: out = 64'b0;
			8'hA0: out = 64'b0;
			8'hA1: out = 64'b0;
			8'hA2: out = 64'b0;
			8'hA3: out = 64'b0;
			8'hA4: out = 64'b0;
			8'hA5: out = 64'b0;
			8'hA6: out = 64'b0;
			8'hA7: out = 64'b0;
			8'hA8: out = 64'b0;
			8'hA9: out = 64'b0;
			8'hAA: out = 64'b0;
			8'hAB: out = 64'b0;
			8'hAC: out = 64'b0;
			8'hAD: out = 64'b0;
			8'hAE: out = 64'b0;
			8'hAF: out = 64'b0;
			8'hB0: out = 64'b0;
			8'hB1: out = 64'b0;
			8'hB2: out = 64'b0;
			8'hB3: out = 64'b0;
			8'hB4: out = 64'b0;
			8'hB5: out = 64'b0;
			8'hB6: out = 64'b0;
			8'hB7: out = 64'b0;
			8'hB8: out = 64'b0;
			8'hB9: out = 64'b0;
			8'hBA: out = 64'b0;
			8'hBB: out = 64'b0;
			8'hBC: out = 64'b0;
			8'hBD: out = 64'b0;
			8'hBE: out = 64'b0;
			8'hBF: out = 64'b0;
			8'hC0: out = 64'b0;
			8'hC1: out = 64'b0;
			8'hC2: out = 64'b0;
			8'hC3: out = 64'b0;
			8'hC4: out = 64'b0;
			8'hC5: out = 64'b0;
			8'hC6: out = 64'b0;
			8'hC7: out = 64'b0;
			8'hC8: out = 64'b0;
			8'hC9: out = 64'b0;
			8'hCA: out = 64'b0;
			8'hCB: out = 64'b0;
			8'hCC: out = 64'b0;
			8'hCD: out = 64'b0;
			8'hCE: out = 64'b0;
			8'hCF: out = 64'b0;
			8'hD0: out = 64'b0;
			8'hD1: out = 64'b0;
			8'hD2: out = 64'b0;
			8'hD3: out = 64'b0;
			8'hD4: out = 64'b0;
			8'hD5: out = 64'b0;
			8'hD6: out = 64'b0;
			8'hD7: out = 64'b0;
			8'hD8: out = 64'b0;
			8'hD9: out = 64'b0;
			8'hDA: out = 64'b0;
			8'hDB: out = 64'b0;
			8'hDC: out = 64'b0;
			8'hDD: out = 64'b0;
			8'hDE: out = 64'b0;
			8'hDF: out = 64'b0;
			8'hE0: out = 64'b0;
			8'hE1: out = 64'b0;
			8'hE2: out = 64'b0;
			8'hE3: out = 64'b0;
			8'hE4: out = 64'b0;
			8'hE5: out = 64'b0;
			8'hE6: out = 64'b0;
			8'hE7: out = 64'b0;
			8'hE8: out = 64'b0;
			8'hE9: out = 64'b0;
			8'hEA: out = 64'b0;
			8'hEB: out = 64'b0;
			8'hEC: out = 64'b0;
			8'hED: out = 64'b0;
			8'hEE: out = 64'b0;
			8'hEF: out = 64'b0;
			8'hF0: out = 64'b0;
			8'hF1: out = 64'b0;
			8'hF2: out = 64'b0;
			8'hF3: out = 64'b0;
			8'hF4: out = 64'b0;
			8'hF5: out = 64'b0;
			8'hF6: out = 64'b0;
			8'hF7: out = 64'b0;
			8'hF8: out = 64'b0;
			8'hF9: out = 64'b0;
			8'hFA: out = 64'b0;
			8'hFB: out = 64'b0;
			8'hFC: out = 64'b0;
			8'hFD: out = 64'b0;
			8'hFE: out = 64'b0;
			8'hFF: out = 64'b0;
			default: out = 64'b0;
		endcase
	end
endmodule
