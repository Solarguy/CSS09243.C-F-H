module rom(out, address);
	output reg [63:0] out;
	input [31:0] address;
	
	always @(address) begin
		if (address[11:0] == 12'hFFF && address[31:20] == 12'h000) begin
			case (address[19:12])
	
	
		// Overclock (Nice!) Test
				0:  out = 32'b11010010100_0000000000000000_01000; // MOVZ X8, 0
				1:  out = 32'b1101001101100000_000000_0100001000; // LSL X8, X8, 0
				2:  out = 32'b11010010100000000000000000100111; // MOVZ X7, 1
				3:  out = 32'b1101001101100000_011000_0011100111; // LSL X7, X7, 24
				4:  out = 32'b11111000000000110000000100000111; // STUR X7, [X8, 48]
				6:  out = 32'b10010100000000000000000000000001; // BL 1
				7:  out = 32'b11010001000001100101011111100000; // SUBI X0, XZR, 405
				8:  out = 32'b11010001000100000000001111100101; // SUBI X5, XZR, 1024
				9:  out = 32'b10110010000001000110011111100010; // ORRI X2, XZR, 281
				10:  out = 32'b10001011000001010000000001000010; // ADD X2, X2, X5
				11:  out = 32'b10001011000001010000000000000000; // ADD X0, X0, X5
				12:  out = 32'b10001011000001010000000010100101; // ADD X5, X5, X5
				13:  out = 32'b10001011000000100000000010100010; // ADD X2, X5, X2
				14:  out = 32'b11010011011000000000010010100101; // LSL X5, X5, 1
				15:  out = 32'b10001011000001010000000000000000; // ADD X0, X0, X5
				16:  out = 32'b11010011011000000000010010100101; // LSL X5, X5, 1
				17:  out = 32'b10001011000001010000000001000010; // ADD X2, X2, X5
				18:  out = 32'b11001011000001010000001111100101; // SUB X5, XZR, X5
				19:  out = 32'b10001011000000100000000000000000; // ADD X0, X0, X2
				20:  out = 32'b10001011000000100000000000000000; // ADD X0, X0, X2
				21:  out = 32'b11111000000000011000000100000000; // STUR X0, [X8, 24]
				22:  out = 32'b11111000000000100000000100000010; // STUR X2, [X8, 32]
				23:  out = 32'b11111000000000101000000100000101; // STUR X5, [X8, 40]
				24:  out = 32'b10010001000000000000001111100000; // ADDI X0, XZR, 0
				25:  out = 32'b10010010000000000000001111100001; // ANDI X1, XZR, 0
				26:  out = 32'b11010010000000000000001111100010; // EORI X2, XZR, 0
				27:  out = 32'b10110010000000000000001111100011; // ORRI X3, XZR, 0
				28:  out = 32'b10101010000111110000001111100100; // ORR X4, X31, X31
				29:  out = 32'b10001010000111110000001111100101; // AND X5, X31, X31
				30:  out = 32'b10001010000111110000001111100110; // AND X6, X31, X31
				31:  out = 32'b11111000010000110000000100000111; // LDUR X7, [X8, 48]
				32:  out = 32'b11010001000000000000010011100111; // SUBI X7, X7, 1
				33:  out = 32'b10110101111111111111111111100111; // CBNZ X7, -1
				34:  out = 32'b11010010100111111111111111100000; // MOVZ X0, 65535
				35:  out = 32'b11010001000000000000011111100001; // SUBI X1, XZR, 1
				36:  out = 32'b11010010100111111111111111100010; // MOVZ X2, 65535
				37:  out = 32'b11010001000000000000011111100011; // SUBI X3, XZR, 1
				38:  out = 32'b11010010100111111111111111100100; // MOVZ X4, 65535
				39:  out = 32'b11010001000000000000011111100101; // SUBI X5, XZR, 1
				40:  out = 32'b11010001000000000000011111100110; // SUBI X6, XZR, 1
				41:  out = 32'b11111000010000110000000100000111; // LDUR X7, [X8, 48]
				42:  out = 32'b11010001000000000000010011100111; // SUBI X7, X7, 1
				43:  out = 32'b10110101111111111111111111100111; // CBNZ X7, -1
				44:  out = 32'b11111000010000011000000100000100; // LDUR X4, [X8, 24]
				45:  out = 32'b11111000010000100000000100000010; // LDUR X2, [X8, 32]
				46:  out = 32'b11111000010000101000000100000101; // LDUR X5, [X8, 40]
				47:  out = 32'b10010001000000000000000001000011; // ADDI X3, X2, 0
				48:  out = 32'b10110010000000010000000001100011; // ORRI X3, X3, 64
				49:  out = 32'b11010010100000000000000100000111; // MOVZ X7, 8
				50:  out = 32'b11001011000001110000000001100011; // SUB X3, X3, X
				51:  out = 32'b11010010100000000000000000100111; // MOVZ X7, 
				52:  out = 32'b11001010000001110000000001100001; // EOR X1, X3, X
				53:  out = 32'b11001011000001010000000000100001; // SUB X1, X1, X5
				54:  out = 32'b10110010000000000000000010000000; // ORRI X0, X4, 0
				55:  out = 32'b11010010100000000000000000000101; // MOVZ X5, 0
				56:  out = 32'b11010010100000000000000000000110; // MOVZ X6, 0
				57:  out = 32'b11111000010000110000000100000111; // LDUR X7, [X8, 48]
				58:  out = 32'b11010001000000000000010011100111; // SUBI X7, X7, 
				59:  out = 32'b10110101111111111111111111100111; // CBNZ X7, -1
				60:  out = 32'b11010110000000000000001111000000; // BR X30

	//input 3 bit number (7) input , compare it with immediate 
	//compare with register that has 1 in it
	
		
		/*
				0: out = 32'b10010001000000000000011101111011; // ADDI X27, X27, 1 				for storing...    movz data in, adjust address LSL,STUR
				1: out = 32'b11010011011000000101001101111011; //LSL X27, X27, 20 
				2: out = 32'b11010010100000000000110001110011; //MOVZ X19, 99    - for 'c'
				3: out = 32'b11111000000000000000001101110011; //STUR X19, [X27, 0]
				4: out = 32'b11010010100000000000111010110100; //MOVZ X20 117		-for 'u'
				5: out = 32'b11010011011000000000011101111011; //LSL X27, X27, 1
				6: out = 32'b11111000000000000000001101110100; //STUR X20, [X27 0]
				7: out = 32'b11010010100000000000111001010011; //MOVZ X19 114		-for 'r'
				8: out = 32'b11010010100000000000000001111011; //MOVZ X27, 3    
				9: out = 32'b11010011011000000101001101111011; //LSL X27 X27, 20
				10: out = 32'b11111000000000000000001101110011; //STUR X19, [X27, 0]
				11: out = 32'b11010010100000000000111001110100; //MOVZ X20, 115 	-for 's'
				12: out = 32'b11010010100000000000000000111011; //MOVZ X27, 1
				13: out = 32'b11010011011000000101101101111011; //LSL X27 X27, 22
				14: out = 32'b11111000000000000000001101110100; //STUR X20 [X27, 0]
				15: out = 32'b11010010100000000000110111110011; //MOVZ X19, 111   - for 'o'
				16: out = 32'b11010010100000000000000010111011; //MOVZ X27 5
				17: out = 32'b11010011011000000101001101111011; //LSL X27 X27, 20
				18: out = 32'b11111000000000000000001101110011; //STUR X19 X27 0
				19: out = 32'b11010010100000000000010000010100; //MOVZ X20 32		-for ' '
				20: out = 32'b11010010100000000000000001111011; //MOVZ X27, 3 
				21: out = 32'b11010011011000000101011101111011; //LSL X27 X27 21
				22: out = 32'b11111000000000000000001101110100; //STUR X20 [X27, 0]
				
				23: out = 32'b11010010100000000000111110010100; //MOVZ X20 124 -for '|'
				24: out = 32'b11010010100000000000000011111011; //MOVZ X27 7
				25: out = 32'b11010011011000000101001101111011; //LSL X27 X27, 20
				26: out = 32'b11111000000000000000001101110100; //STUR X20 [X27, 0];	
				
				27: out = 32'b11010010100000000000110011110011; //MOVZ X19 103 	-for 'g'
				28: out = 32'b11010010100000000000000000111011; //MOVZ X27, 1;
				29: out = 32'b11010011011000000101111101111011; //LSL X27 X27 23
				30: out = 32'b11111000000000000000001101110011; //STUR X19 X27 0
				
				31: out = 32'b11010010100000000000110000110100; //MOVZ X20 97	 	-for 'a'
				32: out = 32'b11010010100000000000000100111011; //MOVZ X27 9
				33: out = 32'b11010011011000000101001101111011; //LSL X27, X27, 20
				34: out = 32'b11111000000000000000001101110100; //STUR X20 [X27, 0];
				
				35: out = 32'b11010010100000000000110111010011; //MOVZ X19 110		-for 'n'
				36: out = 32'b11010010100000000000000101011011; //MOVZ X27 10
				37: out = 32'b11010011011000000101001101111011; //LSL X27, X27, 20 
				38: out = 32'b11111000000000000000001101110011; //STUR X19 X27 0
				
				39: out = 32'b11010010100000000000110010010100; //MOVZ X20 100		-for 'd'
				40: out = 32'b11010010100000000000000101111011; //MOVZ X27 11
				41: out = 32'b11010011011000000101001101111011; //LSL X27, X27, 20 
				42: out = 32'b11111000000000000000001101110100; //STUR X20 [X27, 0];
				
				43: out = 32'b11010010100000000000110110110011; //MOVZ X19 109		-for 'm'
				44: out = 32'b11010010100000000000000110011011; //MOVZ X27 12
				45: out = 32'b11010011011000000101001101111011; //LSL X27, X27, 20 
				46: out = 32'b11111000000000000000001101110011; //STUR X19 X27 0
				
				//Load Registers Recursively in Cookie Clicker Program
				47: out = 32'b11010010100000000000000110010001; //MOVZ X17 12
				48: out = 32'b11010010100000000000000110111011; //MOVZ X27 13
				49: out = 32'b11010011011000000101001101111011; //LSL X27, X27, 20 
				50: out = 32'b11111000000000000000001101110001; //STUR X17 X27 0
			
				51: out = 32'b11010010100000000000000000110010; //MOVZ X18 1
				52: out = 32'b11010010100000000000000111011011; //MOVZ X27 14
				53: out = 32'b11010011011000000101001101111011; //LSL X27, X27, 20 
				54: out = 32'b11111000000000000000001101110010; //STUR X18 X27 0
				
				
				*/
				
				
				
				
				
			/*
				0: out = 32'b10010001000000000011110000000000; // ADDI X0, X0, 15
				1: out = 32'b10010001000000000111110000100001; // ADDI X1, X1, 31
				2: out = 32'b10010001000000000011110001000010; //ADDI X2, X2, 15
				3: out = 32'b11010010100000000000000000100011; //MOVZ X3, 1
				4: out = 32'b11010010100000000000000001000100; //MOVZ X4, 2
				5: out = 32'b10010001000000000000110010100101; // ADDI X5, X5, 3
				6: out = 32'b10010001000000000001000011000110; //ADDI X6, X6, 4
				7: out = 32'b11010010100000000000000010100111; //MOVZ, X7, 5 
				
				*/
				
				
				
			
		/*
				0: out = 32'b10010001000000000011110000000000; // ADDI X0, X0, 15
				1: out = 32'b10010001000000000111110000100001; // ADDI X1, X1, 31
				2: out = 32'b10010001000000000011110001000010; //ADDI X2, X2, 15
				3: out = 32'b10101010001000010000000001000011 ; //ORN X3, X1, X0
				4: out = 32'b11110010000000000011110000011111; // TSTI X31, X0, 15
				5: out = 32'b11101010000000010000000000011111; // TSTR X31, X0, X1
				6: out = 32'b11101011000000010000000000011111; // CMPR X31, X0, X1
				7: out = 32'b11101011000000000000000000111111; // CMPR X31, X1, X0
				8: out = 32'b10010001000000000011000010100101; //ADDI X5, X5, 12
				9: out = 32'b10101010001001010000000001000100; //ORN X4, X5, X2
				10: out = 32'b10010001000000000111110011100111; //ADDI X7, X7, 31
				11: out = 32'b11101011000001110000000000111111; // CMPR  X31, X1, X7
				
*/
			
			/*
			
				// Overclock (Nice!) Test
				// use X8 as the base address of RAM (default is 0x00000000)
				// For example if RAM is at 0x80000000 then change the following two instructions to:
				// MOVZ X8, 8 (put 8 in X8)
				// LSL X8, X8, 28 (shift it 28 times to get 0x80000000)
				0:  out = 32'b11010010100_0000000000000000_01000; // MOVZ X8, 0
				1:  out = 32'b1101001101100000_000000_0100001000; // LSL X8, X8, 0
				// use X11 as the base address of ROM (default is 0x00008000)
				2:  out = 32'b11010010100_0000000000001000_01011; // MOVZ X11, 8
				3:  out = 32'b11010011011000000011000101101011; // LSL X11, X11, 12
				// X7 will hold the delay amount                                        POSSIBLE ISSUE HERE
				4:  out = 32'b11010010100000000000000000100111; // MOVZ X7, 1
				// change the shift amount to change the delay
				// if using a testbench to debug then change the shift amount to 1
				5:  out = 32'b1101001101100000_011000_0011100111; // LSL X7, X7, 24
				6:  out = 32'b11111000000000110000000100000111; // STUR X7, [X8, 48]
				7:  out = 32'b11010001000001100101011111100000; // SUBI X0, XZR, 405
				8:  out = 32'b11010001000100000000001111100101; // SUBI X5, XZR, 1024
				9:  out = 32'b10110010000001000110011111100010; // ORRI X2, XZR, 281
				10:  out = 32'b10001011000001010000000001000010; // ADD X2, X2, X5
				11:  out = 32'b10001011000001010000000000000000; // ADD X0, X0, X5
				12:  out = 32'b10001011000001010000000010100101; // ADD X5, X5, X5
				13:  out = 32'b10001011000000100000000010100010; // ADD X2, X5, X2
				14:  out = 32'b11010011011000000000010010100101; // LSL X5, X5, 1
				15:  out = 32'b10001011000001010000000000000000; // ADD X0, X0, X5
				16:  out = 32'b11010011011000000000010010100101; // LSL X5, X5, 1
				17:  out = 32'b10001011000001010000000001000010; // ADD X2, X2, X5
				18:  out = 32'b11001011000001010000001111100101; // SUB X5, XZR, X5
				19:  out = 32'b10001011000000100000000000000000; // ADD X0, X0, X2
				20:  out = 32'b10001011000000100000000000000000; // ADD X0, X0, X2
				21:  out = 32'b11111000000000011000000100000000; // STUR X0, [X8, 24]
				22:  out = 32'b11111000000000100000000100000010; // STUR X2, [X8, 32]
				23:  out = 32'b11111000000000101000000100000101; // STUR X5, [X8, 40]
				24:  out = 32'b10010001000000000000001111100000; // ADDI X0, XZR, 0
				25:  out = 32'b10010010000000000000001111100001; // ANDI X1, XZR, 0
				26:  out = 32'b11010010000000000000001111100010; // EORI X2, XZR, 0
				27:  out = 32'b10110010000000000000001111100011; // ORRI X3, XZR, 0
				28:  out = 32'b10101010000111110000001111100100; // ORR X4, X31, X31
				29:  out = 32'b10001010000111110000001111100101; // AND X5, X31, X31
				30:  out = 32'b10001010000111110000001111100110; // AND X6, X31, X31
				31:  out = 32'b11111000010000110000000100000111; // LDUR X7, [X8, 48]
				32:  out = 32'b11010001000000000000010011100111; // SUBI X7, X7, 1
			  // 33:  out = 32'b10110101111111111111111110100111; // CBNZ X7, -3
				34:  out = 32'b11010010100111111111111111100000; // MOVZ X0, 65535
				35:  out = 32'b11010001000000000000011111100001; // SUBI X1, XZR, 1
				36:  out = 32'b11010010100111111111111111100010; // MOVZ X2, 65535
				37:  out = 32'b11010001000000000000011111100011; // SUBI X3, XZR, 1
				38:  out = 32'b11010010100111111111111111100100; // MOVZ X4, 65535
				39:  out = 32'b11010001000000000000011111100101; // SUBI X5, XZR, 1
				40:  out = 32'b11010001000000000000011111100110; // SUBI X6, XZR, 1
				41:  out = 32'b11111000010000110000000100000111; // LDUR X7, [X8, 48]
				42:  out = 32'b11010001000000000000010011100111; // SUBI X7, X7, 1
			//	43:  out = 32'b10110101111111111111111110100111; // CBNZ X7, -3
				44:  out = 32'b11111000010000011000000100000100; // LDUR X4, [X8, 24]
				45:  out = 32'b11111000010000100000000100000010; // LDUR X2, [X8, 32]
				46:  out = 32'b11111000010000101000000100000101; // LDUR X5, [X8, 40]
				47:  out = 32'b10010001000000000000000001000011; // ADDI X3, X2, 0
				48:  out = 32'b10110010000000010000000001100011; // ORRI X3, X3, 64
				49:  out = 32'b11010010100000000000000100000111; // MOVZ X7, 8
				50:  out = 32'b11001011000001110000000001100011; // SUB X3, X3, X
				51:  out = 32'b11010010100000000000000000100111; // MOVZ X7, 
				52:  out = 32'b11001010000001110000000001100001; // EOR X1, X3, X
				53:  out = 32'b11001011000001010000000000100001; // SUB X1, X1, X5
				54:  out = 32'b10110010000000000000000010000000; // ORRI X0, X4, 0
				55:  out = 32'b11010010100000000000000000000101; // MOVZ X5, 0
				56:  out = 32'b11010010100000000000000000000110; // MOVZ X6, 0
				57:  out = 32'b11111000010000110000000100000111; // LDUR X7, [X8, 48]
				58:  out = 32'b11010001000000000000010011100111; // SUBI X7, X7, 
				//59:  out = 32'b10110101111111111111111110100111; // CBNZ X7, -3               maybe try -3
				60:  out = 32'b11010110000000000000000101100000; // BR X11
				
				//end overclock tst
		
				
				
				*/
				
				
				
				
				
				
				
				/*0: out = 32'b10010100000000000000000000000011; // BL 3
				1: out = 32'b10010001000000000000010000000000; // ADDI X0, X0, 1
				2: out = 32'b00010111111111111111111111111111; // B -1
				3: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
				4: out = 32'b11010110000000000000001111000000; // BR 30*/
				
				/*0: out = 32'b11010010100000000000000000100001; // MOVZ X1, 1
				1: out = 32'b11010010100000000000000001000010; // MOVZ X2, 2
				2: out = 32'b10001011000000100000000000100100; // ADD X4, X1, X2
				3: out = 32'b11111000000000010000001111100100; // STUR X4, [XZR, 16]
				//5: out = 32'b11111000010000010000001111100101; // LDUR X5, [XZR, 16]
				4: out = 32'b10010100000000000000000000001010; // BL 10
				5: out = 32'b10110101000000000000000000100010; // CBNZ X2, 1
				6: out = 32'b00010100000000000000000000000001; // B 1
				7: out = 32'b00010111111111111111111111111001; // B -7
				8: out = 32'b10110100000000000000000001100001; // CBZ X1, 3
				9: out = 32'b11101011000000100000000000111111; // SUBS XZR, X1, X2
				10: out = 32'b01010100000000000000000000100011; // B.LO 1
				11: out = 32'b11111000000000001000001111100001; // STUR X1, [XZR, 8]
				12: out = 32'b11111000010000001000001111100110; // LDUR X6, [XZR, 8]
				13: out = 32'b11010010000000000000010011100111; // EORI X7, X7, 1
				14: out = 32'b00010111111111111111111111111110; // B -2
				15: out = 32'b10010001000000000000100000100001; // ADDI X1, X1, 2
				16: out = 32'b11010001000000000000010001000010; // SUBI X2, X2, 1
				17: out = 32'b11010110000000000000001111000000; // BR X30*/
				
				/*0: out = 32'b10010001000000000000010000000000; // ADDI X0, X0, 1
				1: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
				2: out = 32'b00010111111111111111111111111111; // B -1*/
				
				/*0: out = 32'b10010001000011111111110000000000; // ADDI X0, X0, 1023
				1: out = 32'b11111000000000000001000000100000; // STUR X0, [X1, 1]
				2: out = 32'b00111000010000000001000000100001; // LDURB X1, [X1, 1]*/
				
				/*0: out = 32'b10010001000000000000110000000000; // ADDI X0, X0, 3
				1: out = 32'b10010001001111111111000000100001; // ADDI X1, X1, -4
				2: out = 32'b10011011000000000000000000100010; // MUL X2, X1, X0*/
				
				/*0: out = 32'b10010001000111111111110000000000; // ADDI X0, X0, 2047
				1: out = 32'b10010001001000000000000000000000; // ADDI X0, X0, 2048
				2: out = 32'b10010001000011111111110000100001; // ADDI X1, X1, 1023
				3: out = 32'b10010001000100000000000000100001; // ADDI X1, X1, 1024
				4: out = 32'b10010001000001111111110001000010; // ADDI X2, X2, 511
				5: out = 32'b10010001000010000000000001000010; // ADDI X2, X2, 512
				6: out = 32'b10010001000000111111110001100011; // ADDI X3, X3, 255
				7: out = 32'b10010001000001000000000001100011; // ADDI X3, X3, 256
				8: out = 32'b10010001000000011111110010000100; // ADDI X4, X4, 127
				9: out = 32'b10010001000000100000000010000100; // ADDI X4, X4, 128
				10: out = 32'b10010001000000001111110010100101; // ADDI X5, X5, 63
				11: out = 32'b10010001000000010000000010100101; // ADDI X5, X5, 64
				12: out = 32'b10010001000000000111110011000110; // ADDI X6, X6, 31
				13: out = 32'b10010001000000001000000011000110; // ADDI X6, X6, 32
				14: out = 32'b10010001000000000011110011100111; // ADDI X7, X7, 15
				15: out = 32'b10010001000000000100000011100111; // ADDI X7, X7, 16
				16: out = 32'b10010001000000000001110100001000; // ADDI X8, X8, 7
				17: out = 32'b10010001000000000010000100001000; // ADDI X8, X8, 8
				18: out = 32'b10010001000000000000110100101001; // ADDI X9, X9, 3
				19: out = 32'b10010001000000000001000100101001; // ADDI X9, X9, 4
				20: out = 32'b10010001000000000000010101001010; // ADDI X10, X10, 1
				21: out = 32'b10010001000000000000100101001010; // ADDI X10, X10, 2
				22: out = 32'b10010001000000000000010101101011; // ADDI X11, X11, 1
				23: out = 32'b10010001001111111111100110001100; // ADDI X12, X12, 4094
				24: out = 32'b10010001001111111111100110001100; // ADDI X12, X12, 4094
				25: out = 32'b10010001000000000000110110001100; // ADDI X12, X12, 3*/
				
				//0: out = 32'b10010001000000000000010000000000; // ADDI X0, X0, 1
				//1: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
				//2: out = 32'b10011010000000010000000000000010; // ADC X2, X0, X1
				//2: out = 32'b10001011000000010000000000000010; // ADD X2, X0, X1
				
				//0: out = 32'b10010001001111111111100001100011;
				//1: out = 32'b11010011011000001101000001100011;
				//2: out = 32'b10010001001111111111100010000100;
				//3: out = 32'b11010011011000001101000010000100;
				//4: out = 32'b10101011000001000000000001100000;
				//0: out = 32'b10010001000000000001000001100011;
				//1: out = 32'b10010001000000000000110010000100;
				//2: out = 32'b11101011000000110000000010000000;
				/*0: out = 32'b10010001001111111111100001100011;
				1: out = 32'b11010011011000000010110001100011;
				2: out = 32'b10010001001111111111100001100011;
				3: out = 32'b11010011011000000010110001100011;
				4: out = 32'b10010001001111111111100001100011;
				5: out = 32'b11010011011000000010110001100011;
				6: out = 32'b10010001001111111111100001100011;
				7: out = 32'b11010011011000000010110001100011;
				8: out = 32'b10010001001111111111100001100011;
				9: out = 32'b11010011011000000010110001100011;
				10: out = 32'b10010001001111111111100001100011;
				11: out = 32'b10010001000000000000010001100011;
				12: out = 32'b10110001000000000000100001100011; // Status checker
				13: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
				14: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1*/
				
				/*0: out = 32'b10010001001111111111110000000000; // ADDI X0, X0, 4095*/
				
				/*0: out = 32'b10010001000000000000010000000000; // ADDI X0, X0, 1
				1: out = 32'b10010100000000000000000000000011; // BL 3
				2: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
				3: out = 32'b00010100000000000000000000000011; // B 3
				4: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
				5: out = 32'b11010110000000000000001111000000; // BR X30
				6: out = 32'b10010001000000000000010001100011; // ADDI X3, X3, 1*/
				
				/*0: out = 32'b10010001000000010001010101001010; // ADDI X10, X10, 69
				1: out = 32'b10110100000000000000000001001001; // CB
				2: out = 32'b10010001000000000000010101101011; // ADDI X11, X11, 1
				3: out = 32'b10010001000000000000010101101011; // ADDI X11, X11, 1
				4: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1*/
				
				/*0: out = 32'b00010100000000000000000000001111; // B 15
				1: out = 32'b10010001000000000000010010100101; // ADDI X5, X5, 1
				2: out = 32'b10010001000000000000011000110001; // ADDI X17, X17, 1
				
				10: out = 32'b10010001000000000000011010010100; // ADDI X20, X20, 1
				11: out = 32'b10010001000000000000011010110101; // ADDI X21, X21, 1
				12: out = 32'b10010001000000000000011011010110; // ADDI X22, X22, 1
				13: out = 32'b10010001000000000000011011110111; // 23
				14: out = 32'b10010001000000000000011100011000; // 24
				15: out = 32'b10010001000000000000011100111001; // 25
				16: out = 32'b10010001000000000000011101011010; // 26
				17: out = 32'b10010001000000000000011101111011;
				18: out = 32'b10010001000000000000011110011100;
				19: out = 32'b10010001000000000000011110111101;
				20: out = 32'b10010001000000000000011111011110;*/
				
				//0: out = 32'b10010001000000000000010000000000; // ADDI X0, X0, 1
				//1: out = 32'b11111000000000000000000000100000; // STUR X1, [X1, 0]
				//2: out = 32'b11111000010000000000000001000010; // LDUR X2, [X2, 0]
				/*0: out = 32'b10010001001010101010101111100000; // ADDI X0, X31, 2730
				1: out = 32'b11010011011000000011000000000000; // LSL X0, X0, 12
				2: out = 32'b10010001001010101010100000000000; // ADDI X0, X0, 2730
				3: out = 32'b11110010100000000000101101000000; // MOVK X0, 90
				4: out = 32'b10010001000000000000010000100001; // ADDI, X1, X1, 1*/
				
				default: out = 32'b10001011000111110000001111111111; // ADD X31, X31, X31
			endcase
		end else begin
			out = 32'bz;
		end
	end
endmodule
