module rom_case(out, address);
	output reg [63:0] out;
	input [31:0] address;
	
	always @(address) begin
		if (address[11:0] == 12'hFFF && address[31:20] == 12'h000) begin
			case (address[19:12])
				0: out = 32'b11010010100000000000000000100001; // MOVZ X1, 1
				1: out = 32'b11010010100000000000000001000010; // MOVZ X2, 2
				2: out = 32'b10001011000000100000000000100100; // ADD X4, X1, X2
				3: out = 32'b11111000000000010000001111100100; // STUR X4, [XZR, 16]
				4: out = 32'b11111000010000010000001111100101; // LDUR X5, [XZR, 16]
				5: out = 32'b10010100000000000000000000001010; // BL 10
				6: out = 32'b10110101000000000000000000100010; // CBNZ X2, 1
				7: out = 32'b00010100000000000000000000000001; // B 1
				8: out = 32'b00010111111111111111111111111001; // B -7
				9: out = 32'b10110100000000000000000001100001; // CBZ X1, 3
				10: out = 32'b11101011000000100000000000111111; // SUBS XZR, X1, X2
				11: out = 32'b01010100000000000000000000100011; // B.LO 1
				12: out = 32'b11111000000000001000001111100001; // STUR X1, [XZR, 8]
				13: out = 32'b11111000010000001000001111100110; // LDUR X6, [XZR, 8]
				14: out = 32'b11010010000000000000010011100111; // EORI X7, X7, 1
				15: out = 32'b00010111111111111111111111111110; // B -2
				16: out = 32'b10010001000000000000100000100001; // ADDI X1, X1, 2
				17: out = 32'b11010001000000000000010001000010; // SUBI X2, X2, 1
				18: out = 32'b11010110000000000000001111000000; // BR X30
				
				/*0: out = 32'b10010001000000000000010000000000; // ADDI X0, X0, 1
				1: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
				2: out = 32'b00010111111111111111111111111111; // B -1*/
				
				/*0: out = 32'b10010001000011111111110000000000; // ADDI X0, X0, 1023
				1: out = 32'b11111000000000000001000000100000; // STUR X0, [X1, 1]
				2: out = 32'b00111000010000000001000000100001; // LDURB X1, [X1, 1]*/
				
				/*0: out = 32'b10010001000000000000110000000000; // ADDI X0, X0, 3
				1: out = 32'b10010001001111111111000000100001; // ADDI X1, X1, -4
				2: out = 32'b10011011000000000000000000100010; // MUL X2, X1, X0*/
				
				/*0: out = 32'b10010001000111111111110000000000; // ADDI X0, X0, 2047
				1: out = 32'b10010001001000000000000000000000; // ADDI X0, X0, 2048
				2: out = 32'b10010001000011111111110000100001; // ADDI X1, X1, 1023
				3: out = 32'b10010001000100000000000000100001; // ADDI X1, X1, 1024
				4: out = 32'b10010001000001111111110001000010; // ADDI X2, X2, 511
				5: out = 32'b10010001000010000000000001000010; // ADDI X2, X2, 512
				6: out = 32'b10010001000000111111110001100011; // ADDI X3, X3, 255
				7: out = 32'b10010001000001000000000001100011; // ADDI X3, X3, 256
				8: out = 32'b10010001000000011111110010000100; // ADDI X4, X4, 127
				9: out = 32'b10010001000000100000000010000100; // ADDI X4, X4, 128
				10: out = 32'b10010001000000001111110010100101; // ADDI X5, X5, 63
				11: out = 32'b10010001000000010000000010100101; // ADDI X5, X5, 64
				12: out = 32'b10010001000000000111110011000110; // ADDI X6, X6, 31
				13: out = 32'b10010001000000001000000011000110; // ADDI X6, X6, 32
				14: out = 32'b10010001000000000011110011100111; // ADDI X7, X7, 15
				15: out = 32'b10010001000000000100000011100111; // ADDI X7, X7, 16
				16: out = 32'b10010001000000000001110100001000; // ADDI X8, X8, 7
				17: out = 32'b10010001000000000010000100001000; // ADDI X8, X8, 8
				18: out = 32'b10010001000000000000110100101001; // ADDI X9, X9, 3
				19: out = 32'b10010001000000000001000100101001; // ADDI X9, X9, 4
				20: out = 32'b10010001000000000000010101001010; // ADDI X10, X10, 1
				21: out = 32'b10010001000000000000100101001010; // ADDI X10, X10, 2
				22: out = 32'b10010001000000000000010101101011; // ADDI X11, X11, 1
				23: out = 32'b10010001001111111111100110001100; // ADDI X12, X12, 4094
				24: out = 32'b10010001001111111111100110001100; // ADDI X12, X12, 4094
				25: out = 32'b10010001000000000000110110001100; // ADDI X12, X12, 3*/
				
				//0: out = 32'b10010001000000000000010000000000; // ADDI X0, X0, 1
				//1: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
				//2: out = 32'b10011010000000010000000000000010; // ADC X2, X0, X1
				//2: out = 32'b10001011000000010000000000000010; // ADD X2, X0, X1
				
				//0: out = 32'b10010001001111111111100001100011;
				//1: out = 32'b11010011011000001101000001100011;
				//2: out = 32'b10010001001111111111100010000100;
				//3: out = 32'b11010011011000001101000010000100;
				//4: out = 32'b10101011000001000000000001100000;
				//0: out = 32'b10010001000000000001000001100011;
				//1: out = 32'b10010001000000000000110010000100;
				//2: out = 32'b11101011000000110000000010000000;
				/*0: out = 32'b10010001001111111111100001100011;
				1: out = 32'b11010011011000000010110001100011;
				2: out = 32'b10010001001111111111100001100011;
				3: out = 32'b11010011011000000010110001100011;
				4: out = 32'b10010001001111111111100001100011;
				5: out = 32'b11010011011000000010110001100011;
				6: out = 32'b10010001001111111111100001100011;
				7: out = 32'b11010011011000000010110001100011;
				8: out = 32'b10010001001111111111100001100011;
				9: out = 32'b11010011011000000010110001100011;
				10: out = 32'b10010001001111111111100001100011;
				11: out = 32'b10010001000000000000010001100011;
				12: out = 32'b10110001000000000000100001100011; // Status checker
				13: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
				14: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1*/
				
				/*0: out = 32'b10010001001111111111110000000000; // ADDI X0, X0, 4095*/
				
				/*0: out = 32'b10010001000000000000010000000000; // ADDI X0, X0, 1
				1: out = 32'b10010100000000000000000000000011; // BL 3
				2: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1
				3: out = 32'b00010100000000000000000000000011; // B 3
				4: out = 32'b10010001000000000000010001000010; // ADDI X2, X2, 1
				5: out = 32'b11010110000000000000001111000000; // BR X30
				6: out = 32'b10010001000000000000010001100011; // ADDI X3, X3, 1*/
				
				/*0: out = 32'b10010001000000010001010101001010; // ADDI X10, X10, 69
				1: out = 32'b10110100000000000000000001001001; // CB
				2: out = 32'b10010001000000000000010101101011; // ADDI X11, X11, 1
				3: out = 32'b10010001000000000000010101101011; // ADDI X11, X11, 1
				4: out = 32'b10010001000000000000010000100001; // ADDI X1, X1, 1*/
				
				/*0: out = 32'b00010100000000000000000000001111; // B 15
				1: out = 32'b10010001000000000000010010100101; // ADDI X5, X5, 1
				2: out = 32'b10010001000000000000011000110001; // ADDI X17, X17, 1
				
				10: out = 32'b10010001000000000000011010010100; // ADDI X20, X20, 1
				11: out = 32'b10010001000000000000011010110101; // ADDI X21, X21, 1
				12: out = 32'b10010001000000000000011011010110; // ADDI X22, X22, 1
				13: out = 32'b10010001000000000000011011110111; // 23
				14: out = 32'b10010001000000000000011100011000; // 24
				15: out = 32'b10010001000000000000011100111001; // 25
				16: out = 32'b10010001000000000000011101011010; // 26
				17: out = 32'b10010001000000000000011101111011;
				18: out = 32'b10010001000000000000011110011100;
				19: out = 32'b10010001000000000000011110111101;
				20: out = 32'b10010001000000000000011111011110;*/
				
				//0: out = 32'b10010001000000000000010000000000; // ADDI X0, X0, 1
				//1: out = 32'b11111000000000000000000000100000; // STUR X1, [X1, 0]
				//2: out = 32'b11111000010000000000000001000010; // LDUR X2, [X2, 0]
				/*0: out = 32'b10010001001010101010101111100000; // ADDI X0, X31, 2730
				1: out = 32'b11010011011000000011000000000000; // LSL X0, X0, 12
				2: out = 32'b10010001001010101010100000000000; // ADDI X0, X0, 2730
				3: out = 32'b11110010100000000000101101000000; // MOVK X0, 90
				4: out = 32'b10010001000000000000010000100001; // ADDI, X1, X1, 1*/
				default: out = 32'b10001011000111110000001111111111; // ADD X31, X31, X31
			endcase
		end else begin
			out = 32'bz;
		end
	end
endmodule
